�<Table name="AlbumCopy" schema="dbo"><PrimaryKey /><Column name="AlbumId" datatype="int" default="" length="0" notnull="1" precision="10" scale="0" auto_increment="0" primary_key="1"><Type datatype="string" length="50" unicode="0" binary="0" varlength="1" /></Column><Column name="Title" datatype="nvarchar" default="" length="160" notnull="1" precision="0" scale="0" auto_increment="0" primary_key="0"><Type datatype="string" length="50" unicode="0" binary="0" varlength="1" /></Column><Column name="ArtistId" datatype="int" default="" length="0" notnull="1" precision="10" scale="0" auto_increment="0" primary_key="0"><Type datatype="string" length="50" unicode="0" binary="0" varlength="1" /></Column></Table>    	%For Those About To Rock We Salute You       	Balls to the Wall       	Restless and Wild       	Let There Be Rock       	Big Ones       	Jagged Little Pill       	Facelift       	Warner 25 Anos    	   	Plays Metallica By Four Cellos    
   	
Audioslave       	Out Of Exile       	BackBeat Soundtrack	       	The Best Of Billy Cobham
       	(Alcohol Fueled Brewtality Live! [Disc 1]       	(Alcohol Fueled Brewtality Live! [Disc 2]       	Black Sabbath       	Black Sabbath Vol. 4 (Remaster)       	
Body Count       	Chemical Wedding       	0The Best Of Buddy Guy - The Millenium Collection       	Prenda Minha       	Sozinho Remix Ao Vivo       	Minha Historia       	Afrociberdelia       	Da Lama Ao Caos       	Acústico MTV [Live]       	Cidade Negra - Hits       	Na Pista       	Axé Bahia 2001       	BBC Sessions [Disc 1] [Live]       	
Bongo Fury        	Carnaval 2001    !   	Chill: Brazil (Disc 1)    "   	Chill: Brazil (Disc 2)    #   	Garage Inc. (Disc 1)2    $   	Greatest Hits II3    %   	Greatest Kiss4    &   	Heart of the Night5    '   	International Superhits6    (   	Into The Light7    )   	Meus Momentos8    *   	Minha História9    +   	"MK III The Final Concerts [Disc 1]:    ,   	Physical Graffiti [Disc 1]    -   	Sambas De Enredo 2001    .   	Supernatural;    /   	The Best of Ed Motta%    0   	"The Essential Miles Davis [Disc 1]D    1   	"The Essential Miles Davis [Disc 2]D    2   	The Final Concerts (Disc 2):    3   	Up An' AtomE    4   	 Vinícius De Moraes - Sem LimiteF    5   	Vozes do MPB    6   	Chronicle, Vol. 1L    7   	Chronicle, Vol. 2L    8   	-Cássia Eller - Coleção Sem Limite [Disc 2]M    9   	#Cássia Eller - Sem Limite [Disc 1]M    :   	Come Taste The Band:    ;   	Deep Purple In Rock:    <   	Fireball:    =   	?Knocking at Your Back Door: The Best Of Deep Purple in the 80's:    >   	Machine Head:    ?   	Purpendicular:    @   	Slaves And Masters:    A   	Stormbringer:    B   	The Battle Rages On:    C   	"Vault: Def Leppard's Greatest HitsN    D   	OutbreakO    E   	Djavan Ao Vivo - Vol. 02P    F   	Djavan Ao Vivo - Vol. 1P    G   	Elis Regina-Minha História)    H   	The Cream Of ClaptonQ    I   		UnpluggedQ    J   	Album Of The YearR    K   	
Angel DustR    L   	"King For A Day Fool For A LifetimeR    M   	The Real ThingR    N   	Deixa EntrarS    O   	In Your Honor [Disc 1]T    P   	In Your Honor [Disc 2]T    Q   	
One By OneT    R   	The Colour And The ShapeT    S   	*My Way: The Best Of Frank Sinatra [Disc 1]U    T   	Roda De FunkV    U   	As Canções de Eu Tu Eles    V   	Quanta Gente Veio Ver (Live)    W   	)Quanta Gente Veio ver--Bônus De Carnaval    X   	FacelessW    Y   	American Idiot6    Z   	Appetite for DestructionX    [   	Use Your Illusion IX    \   	Use Your Illusion IIX    ]   	
Blue MoodsY    ^   	A Matter of Life and DeathZ    _   	A Real Dead OneZ    `   	A Real Live OneZ    a   	Brave New WorldZ    b   	Dance Of DeathZ    c   	Fear Of The DarkZ    d   	Iron MaidenZ    e   	KillersZ    f   	Live After DeathZ    g   	Live At Donington 1992 (Disc 1)Z    h   	Live At Donington 1992 (Disc 2)Z    i   	No Prayer For The DyingZ    j   	Piece Of MindZ    k   	
PowerslaveZ    l   	Rock In Rio [CD1]Z    m   	Rock In Rio [CD2]Z    n   	Seventh Son of a Seventh SonZ    o   	Somewhere in TimeZ    p   	The Number of The BeastZ    q   	The X FactorZ    r   	
Virtual XIZ    s   	Sex Machine[    t   	Emergency On Planet Earth\    u   	Synkronized\    v   	The Return Of The Space Cowboy\    w   	Get Born]    x   	Are You Experienced?^    y   	#Surfing with the Alien (Remastered)_    z   	Jorge Ben Jor 25 Anos.    {   	Jota Quest-1995`    |   		Cafezinhoa    }   	Living After Midnightb    ~   	Unplugged [Live]4       	BBC Sessions [Disc 2] [Live]    �   	Coda    �   	Houses Of The Holy    �   	In Through The Out Door    �   	IV    �   	Led Zeppelin I    �   	Led Zeppelin II    �   	Led Zeppelin III    �   	Physical Graffiti [Disc 2]    �   	Presence    �   	"The Song Remains The Same (Disc 1)    �   	"The Song Remains The Same (Disc 2)    �   	*A TempestadeTempestade Ou O Livro Dos Diasc    �   	Mais Do Mesmoc    �   	Greatest Hitsd    �   	1Lulu Santos - RCA 100 Anos De Música - Álbum 01e    �   	1Lulu Santos - RCA 100 Anos De Música - Álbum 02e    �   	Misplaced Childhoodf    �   	Barulhinho Bomg    �   	1Seek And Shall Find: More Of The Best (1963-1981)h    �   	The Best Of Men At Worki    �   	Black Album2    �   	Garage Inc. (Disc 2)2    �   	Kill 'Em All2    �   	Load2    �   	Master Of Puppets2    �   	ReLoad2    �   	Ride The Lightning2    �   		St. Anger2    �   	...And Justice For All2    �   	Miles AheadD    �   	Milton Nascimento Ao Vivo*    �   	Minas*    �   	Ace Of Spadesj    �   	
Demorou...l    �   	Motley Crue Greatest Hitsm    �   	*From The Muddy Banks Of The Wishkah [Live]n    �   		Nevermindn    �   	Compositoreso    �   	Olodump    �   	Acústico MTVq    �   	
Arquivo IIq    �   	Arquivo Os Paralamas Do Sucessoq    �   	Bark at the Moon (Remastered)r    �   	Blizzard of Ozzr    �   	Diary of a Madman (Remastered)r    �   	No More Tears (Remastered)r    �   	Tributer    �   	Walking Into Clarksdales    �   	Original Soundtracks 1t    �   	The Beast Liveu    �   	Live On Two Legs [Live]v    �   		Pearl Jamv    �   	Riot Actv    �   	Tenv    �   	Vs.v    �   	Dark Side Of The Moonx    �   	)Os Cães Ladram Mas A Caravana Não Páray    �   	Greatest Hits I3    �   	News Of The World3    �   	Out Of Timez    �   	Green|    �   	New Adventures In Hi-Fi|    �   	!The Best Of R.E.M.: The IRS Years|    �   	Cesta Básica}    �   	Raul Seixas~    �   	Blood Sugar Sex Magik    �   	
By The Way    �   	Californication    �   	Retrospective I (1974-1980)�    �   	Santana - As Years Go By;    �   	Santana Live;    �   	Maquinarama�    �   	O Samba Poconé�    �   	Judas 0: B-Sides and Rarities�    �   	Rotten Apples: Greatest Hits�    �   	A-Sides�    �   	Morning Dance5    �   	In Step�    �   	Core�    �   		Mezmerize�    �   	[1997] Black Light Syndrome�    �   	Live [Disc 1]�    �   	Live [Disc 2]�    �   	The Singles�    �   	Beyond Good And Evil�    �   	LPure Cult: The Best Of The Cult (For Rockers, Ravers, Lovers & Sinners) [UK]�    �   		The Doors�    �   	The Police Greatest Hits�    �   	Hot Rocks, 1964-1971 (Disc 1)�    �   	No Security�    �   	Voodoo Lounge�    �   	Tangents�    �   	Transmission�    �   	(My Generation - The Very Best Of The Who�    �   	Serie Sem Limite (Disc 1)�    �   	Serie Sem Limite (Disc 2)�    �   		Acústico�    �   	Volume Dois�    �   	&Battlestar Galactica: The Story So Far�    �   	Battlestar Galactica, Season 3�    �   	Heroes, Season 1�    �   	Lost, Season 3�    �   	Lost, Season 1�    �   	Lost, Season 2�    �   	Achtung Baby�    �   	All That You Can't Leave Behind�    �   	B-Sides 1980-1990�    �   	How To Dismantle An Atomic Bomb�    �   	Pop�    �   	Rattle And Hum�    �   	The Best Of 1980-1990�    �   	War�    �   	Zooropa�    �   	"UB40 The Best Of - Volume Two [UK]�    �   	
Diver Down�    �   	The Best Of Van Halen, Vol. I�    �   		Van Halen�    �   	Van Halen III�    �   	
Contraband�    �   	Vinicius De MoraesH    �   	Ao Vivo [IMPORT]�    �   	The Office, Season 1�    �   	The Office, Season 2�    �   	The Office, Season 3�    �   		Un-Led-Ed�    �   	(Battlestar Galactica (Classic), Season 1�    �   	Aquaman�    �   	@Instant Karma: The Amnesty International Campaign to Save Darfur�       	Speak of the Devilr      	G20th Century Masters - The Millennium Collection: The Best of Scorpions�      	House of Pain�      	DRadio Brasil (O Som da Jovem Vanguarda) - Seleccao de Henrique Amaro$      	Cake: B-Sides and Rarities�      	LOST, Season 4�      	Quiet Songs�      	Muso Ko�      	Realize�    	  	Every Kind of Light�    
  	Duos II�      	Worlds�      	The Best of Beethoven�      	Temple of the Dog�      	Carry On�      	Revelations      	9Adorate Deum: Gregorian Chant from the Proper of the Mass�      	Allegri: Miserere�      	Pachelbel: Canon & Gigue�      	Vivaldi: The Four Seasons�      	Bach: Violin Concertos�      	Bach: Goldberg Variations�      	Bach: The Cello Suites�      	 Handel: The Messiah (Highlights)�      	!The World of Classical Favourites�      	#Sir Neville Marriner: A Celebration�      	Mozart: Wind Concertos�      	Haydn: Symphonies 99 - 104�      	Beethoven: Symhonies Nos. 5 & 6�      	A Soprano Inspired�      	Great Opera Choruses�      	Wagner: Favourite Overtures�       	'Fauré: Requiem, Ravel: Pavane & Others�    !  	Tchaikovsky: The Nutcracker�    "  	The Last Night of the Proms�    #  	&Puccini: Madama Butterfly - Highlights�    $  	8Holst: The Planets, Op. 32 & Vaughan Williams: Fantasies�    %  	Pavarotti's Opera Made Easy�    &  	MGreat Performances - Barber's Adagio and Other Romantic Favorites for Strings�    '  	Carmina Burana�    (  	A Copland Celebration, Vol. I�    )  	 Bach: Toccata & Fugue in D Minor�    *  	Prokofiev: Symphony No.1�    +  	Scheherazade�    ,  	Bach: The Brandenburg Concertos�    -  	"Chopin: Piano Concertos Nos. 1 & 2�    .  	Mascagni: Cavalleria Rusticana�    /  	Sibelius: Finlandia�    0  	.Beethoven Piano Sonatas: Moonlight & Pastorale�    1  	?Great Recordings of the Century - Mahler: Das Lied von der Erde�    2  	3Elgar: Cello Concerto & Vaughan Williams: Fantasias�    3  	 Adams, John: The Chairman Dances�    4  	_Tchaikovsky: 1812 Festival Overture, Op.49, Capriccio Italien & Beethoven: Wellington's Victory�    5  	4Palestrina: Missa Papae Marcelli & Allegri: Miserere�    6  	Prokofiev: Romeo & Juliet�    7  	Strauss: Waltzes�    8  	Berlioz: Symphonie Fantastique�    9  	Bizet: Carmen Highlights�    :  	English Renaissance�    ;  	=Handel: Music for the Royal Fireworks (Original Version 1749)�    <  	:Grieg: Peer Gynt Suites & Sibelius: Pelléas et Mélisande�    =  	Mozart Gala: Famous Arias�    >  	SCRIABIN: Vers la flamme�    ?  	2Armada: Music from the Courts of England and Spain�    @  	Mozart: Symphonies Nos. 40 & 41�    A  	Back to Black�    B  	Frank�    C  	%Carried to Dust (Bonus Track Version)�    D  	)Beethoven: Symphony No. 6 'Pastoral' Etc.�    E  	 Bartok: Violin & Viola Concertos�    F  	&Mendelssohn: A Midsummer Night's Dream    G  	"Bach: Orchestral Suites Nos. 1 - 4   H  	-Charpentier: Divertissements, Airs & Concerts   I  	South American Getaway   J  	Górecki: Symphony No. 3   K  	Purcell: The Fairy Queen   L  	The Ultimate Relexation Album   M  	!Purcell: Music for the Queen Mary   N  	Weill: The Seven Deadly Sins   O  	VJ.S. Bach: Chaconne, Suite in E Minor, Partita in E Major & Prelude, Fugue and Allegro	   P  	<Prokofiev: Symphony No.5 & Stravinksy: Le Sacre Du Printemps�    Q  	 Szymanowski: Piano Works, Vol. 1
   R  	Nielsen: The Six Symphonies   S  	7Great Recordings of the Century: Paganini's 24 Caprices   T  	,Liszt - 12 Études D'Execution Transcendante   U  	CGreat Recordings of the Century - Shubert: Schwanengesang, 4 Lieder   V  	=Locatelli: Concertos for Violin, Strings and Continuo, Vol. 3   W  	Respighi:Pines of Rome�    X  	<Schubert: The Late String Quartets & String Quintet (3 CD's)   Y  	Monteverdi: L'Orfeo   Z  	Mozart: Chamber Music   [  	2Koyaanisqatsi (Soundtrack from the Motion Picture)  